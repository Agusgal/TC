C:\Users\Msrt\Documents\GitHub\TC\TP3\Ej3\Simulaciones\SapWin\ampIns.sch
R3 5 1 1
R4 1 3 1
R6 3 2 1
R7 2 6 1
EO1 5 0 1 10 1e6
EO2 6 0 2 11 1e6
R5 3 4 1
EO4 4 0 0 7 1e6
R1 8 5 1
R2 12 8 1
R8 9 6 1
R9 7 9 1
EO3 12 0 8 9 1e6
V1 10 0 AC 1
V2 11 0 AC 1
.AC DEC 100 1 1000
.PROBE
.END
